** Profile: "SCHEMATIC1-varsen"  [ d:\anul 2.2\sem 2\cad\proiect\proiectfinal-pspicefiles\schematic1\varsen.sim ] 

** Creating circuit file "varsen.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../proiectfinal-pspicefiles/redled.lib" 
* From [PSPICE NETLIST] section of C:\Users\stefa\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\22.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10m 0 
.STEP LIN PARAM r 50k 60k 1k 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
